// DE1_SoC_QSYS.v

// Generated using ACDS version 15.0 145

`timescale 1 ps / 1 ps
module DE1_SoC_QSYS (
		input   wire       clk_clk,                        //Original Reforence clock:50MHz
		input   wire       reset_reset_n,                  //reset signal for whole system: KEY0  
		input   wire [9:0] sw_external_connection_export,  //10 FPGA switches--RESERVED NOW
		input   wire [2:0] sw_ADC_pin_select,
		
		output  wire       pll_sys_locked_export,          //pll_sys_locked.export  ???Just keep it
		
		//--------------------ADC----------------------------------------------------
		input   wire       adc_reset_n,
		output  wire[11:0] ADCout,
		
		output  wire       wait_measure_done,
		output  wire       pll_sys_outclk1_clk,  //40MHz
		
		output  wire       adc_ltc2308_conduit_end_CONVST, // adc_ltc2308_conduit_end.CONVST
		output  wire       adc_ltc2308_conduit_end_SCK,    //                        .SCK
		output  wire       adc_ltc2308_conduit_end_SDI,    //                        .SDI
		input   wire       adc_ltc2308_conduit_end_SDO,    //                        .SDO
		
		//-------------------SDRAM---------------------------------------------------------
		output wire       pll_sys_outclk0_clk,             //100MHz clock for SDRAM
		
		//-------------------SDRAM---------------------------------------------------------
		output wire       pll_sys_outclk2_clk              //25MHz clock for VGA display
	);

	//wire    pll_sys_outclk0_clk;            // pll_sys:outclk_0 -> [adc_ltc2308:slave_clk, rst_controller:clk, sw:clk, sysid_qsys:clock]
	//wire    pll_sys_outclk1_clk;            // pll_sys:outclk_1 -> adc_ltc2308:adc_clk
	wire    rst_controller_reset_out_reset; // rst_controller:reset_out -> [adc_ltc2308:slave_reset_n, sw:reset_n, sysid_qsys:reset_n]

	adc_ltc2308_fifo adc_ltc2308 (
		.slave_chipselect_n (),                                //          slave.chipselect_n
		.slave_read_n       (),                                //               .read_n
		.slave_readdata     (),                                //               .readdata
		.slave_addr         (),                                //               .address
		.slave_wrtie_n      (),                                //               .write_n
		.slave_wriredata    (),                                //               .writedata
		.ADC_CONVST         (adc_ltc2308_conduit_end_CONVST),  //    conduit_end.export
		.ADC_SCK            (adc_ltc2308_conduit_end_SCK),     //               .export
		.ADC_SDI            (adc_ltc2308_conduit_end_SDI),     //               .export
		.ADC_SDO            (adc_ltc2308_conduit_end_SDO),     //               .export
		.slave_reset_n      (~rst_controller_reset_out_reset), //     reset_sink.reset_n
		.slave_clk          (pll_sys_outclk0_clk),             //     clock_sink.clk
		.adc_clk            (pll_sys_outclk1_clk),             // clock_sink_adc.clk
		
		//===============Added for ADC values==========================================
		.sw_ADC_pin_select  (sw_ADC_pin_select),
		.ADCout             (ADCout),
		.adc_reset_n        (adc_reset_n),
		.wait_measure_done  (wait_measure_done)
	);

	DE1_SoC_QSYS_pll_sys pll_sys (
		.refclk   (clk_clk),               //  refclk.clk
		.rst      (~reset_reset_n),        //   reset.reset
		.outclk_0 (pll_sys_outclk0_clk),   // outclk0.clk  100MHz
		.outclk_1 (pll_sys_outclk1_clk),   // outclk1.clk  40MHz
		.outclk_2 (pll_sys_outclk2_clk),   // outclk2.clk  25MHz   ???suspicious
		.locked   (pll_sys_locked_export)  //  locked.export
	);

	DE1_SoC_QSYS_sw sw (
		.clk        (pll_sys_outclk0_clk),             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset), //               reset.reset_n
		.address    (),                                //                  s1.address
		.write_n    (),                                //                    .write_n
		.writedata  (),                                //                    .writedata
		.chipselect (),                                //                    .chipselect
		.readdata   (),                                //                    .readdata
		.in_port    (sw_external_connection_export),   // external_connection.export
		.irq        ()                                 //                 irq.irq
	);

	DE1_SoC_QSYS_sysid_qsys sysid_qsys (
		.clock    (pll_sys_outclk0_clk),             //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset), //         reset.reset_n
		.readdata (),                                // control_slave.readdata
		.address  ()                                 //              .address
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (pll_sys_outclk0_clk),            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
